`ifndef _global_vh_
`define _global_vh_

/**** Memory setup ****/
`define MEM_SIZE     'h10_0000

`define CHANNEL_SIZE    8
`define PIXEL_SIZE      8

/**** Input/output files ****/
`define IFILE       "imgs/stackable.bmp"
`define OFILE       "out/stackable17.bmp"

/**** Testbench setup ****/
`define SIM_TIME 2_000_000

`endif
